`include "parameter.v"
// fpga4student.com 
// FPGA projects, VHDL projects, Verilog projects 
// Verilog code for RISC Processor 
// Verilog code for Instruction Memory
module Instruction_Memory(
  input[7:0] pc,
 output[15:0] instruction
);

 reg [`col - 1:0] memory [`row_i - 1:0];
  wire [7 : 0] rom_addr = pc;
 initial
 begin
  $readmemb("test.prog", memory,0,14);
 end
 assign instruction =  memory[rom_addr]; 

endmodule